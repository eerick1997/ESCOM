module contdec ( 
	clr,
	clk,
	f,
	c,
	display
	) ;

input  clr;
input  clk;
input [3:0] f;
inout [2:0] c;
inout [6:0] display;
