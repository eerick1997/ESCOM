module ffrs ( 
	r,
	s,
	clk,
	pre,
	clr,
	q,
	nq
	) ;

input  r;
input  s;
input  clk;
input  pre;
input  clr;
inout  q;
inout  nq;
