module allff ( 
	clk,
	clr,
	control,
	q
	) ;

input  clk;
input  clr;
input  control;
inout [7:0] q;
