library ieee;
use ieee.std_logic_1164.all;

entity codec is port(
	clk, clr: in std_logic;
	--ent: in std_logic_vector (1 downto 0);

	--Entrada para cargar dato
	carga: in std_logic_vector (3 downto 0);

	y: in std_logic_vector (1 downto 0);
	display: inout std_logic_vector (6 downto 0)
);
end entity;

architecture a_codec of codec is 
constant dig0: std_logic_vector (6 downto 0):= "0000001";
constant dig1: std_logic_vector (6 downto 0):= "1001111";
constant dig2: std_logic_vector (6 downto 0):= "0010101";
constant dig3: std_logic_vector (6 downto 0):= "0000110";
constant dig4: std_logic_vector (6 downto 0):= "1001100";
constant dig5: std_logic_vector (6 downto 0):= "0100100";
constant dig6: std_logic_vector (6 downto 0):= "0100000";
constant dig7: std_logic_vector (6 downto 0):= "0001111";
constant dig8: std_logic_vector (6 downto 0):= "0000000";
constant dig9: std_logic_vector (6 downto 0):= "0001100";
begin
	process(clk,clr,y,display) begin
		if(clr = '0') then
			display <= dig0;
		elsif(clk'event and clk = '1') then
			case y is
				when "00" => display <= display;
				when "01" => 
					case display is
						when dig0 => display <= dig1;
						when dig1 => display <= dig2;
						when dig2 => display <= dig3;
						when dig3 => display <= dig4;
						when dig4 => display <= dig5;
						when dig5 => display <= dig6;
						when dig6 => display <= dig7;
						when dig7 => display <= dig8;
						when dig8 => display <= dig9;
						when dig9 => display <= dig0;
						when others => display <= dig0;
					end case;
				when "10" =>
					case display is
						when dig0 => display <= dig9;
						when dig9 => display <= dig8;
  					    when dig8 => display <= dig7;
						when dig7 => display <= dig6;
						when dig6 => display <= dig5;
						when dig5 => display <= dig4;
						when dig4 => display <= dig3;
						when dig3 => display <= dig2;
						when dig2 => display <= dig1;
						when dig1 => display <= dig0;
						when others => display <= dig0;
					end case;

				 when others =>
				 	--Decodificador BCD 7 seg
					case carga is
						when "0000" => display <= dig0;--State A
						when "0001" => display <= dig1;--State B
						when "0010" => display <= dig2;--State C
						when "0011" => display <= dig3;--State D
						when "0100" => display <= dig4;--State E
						when "0101" => display <= dig5;--State F
						when "0110" => display <= dig6;--State G
						when "0111" => display <= dig7;--State H
						when "1000" => display <= dig8;--State I
						when "1001" => display <= dig9;--State J
						when others => display <= dig0;
					end case;
			end case;
		end if;
	end process;
end a_codec;
