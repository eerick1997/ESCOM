module registros ( 
	a,
	b,
	c,
	sa,
	sb,
	clk,
	clr,
	control
	) ;

inout [3:0] a;
inout [3:0] b;
inout  c;
inout  sa;
inout  sb;
input  clk;
input  clr;
input  control;
