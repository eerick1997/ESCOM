module fft ( 
	t,
	clk,
	pre,
	clr,
	q,
	nq
	) ;

input  t;
input  clk;
input  pre;
input  clr;
inout  q;
inout  nq;
