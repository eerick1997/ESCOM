module contdec ( 
	clr,
	clk,
	control,
	display
	) ;

input  clr;
input  clk;
input  control;
inout [6:0] display;
