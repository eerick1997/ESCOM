library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity PILA is
	GENERIC(
		BITS: INTEGER := 16;
		ADDR: INTEGER := 4
	);
	
	PORT(
		CLK, CLR: IN STD_LOGIC;
		WPC, UP, DW: IN STD_LOGIC;
		D: IN STD_LOGIC_VECTOR(BITS-1 DOWNTO 0);
		STACK_POINTER: INOUT STD_LOGIC_VECTOR(ADDR-1 DOWNTO 0);
		Q: INOUT STD_LOGIC_VECTOR(BITS-1 DOWNTO 0)
	);
end PILA;

architecture PROGRAMA of PILA is
TYPE MEMORY IS ARRAY (0 TO 2**ADDR-1) OF STD_LOGIC_VECTOR(D'RANGE);
SIGNAL STACKS: MEMORY;
SIGNAL DOUT: STD_LOGIC_VECTOR(BITS-1 DOWNTO 0);
begin
	PSP: PROCESS(CLK, CLR) BEGIN
		IF(CLR = '1') THEN
			STACK_POINTER <= (OTHERS => '0');
		ELSIF (RISING_EDGE(CLK)) THEN
			IF(UP = '1') THEN
				STACK_POINTER <= STACK_POINTER + 1;
			ELSIF(DW = '1') THEN
				STACK_POINTER <= STACK_POINTER - 1;
			END IF;
		END IF;
	END PROCESS PSP;

	PPC: PROCESS(CLK, CLR) BEGIN
		IF(CLR = '1') THEN
			Q <= (OTHERS => '0');
		ELSIF(RISING_EDGE(CLK)) THEN
			IF(WPC = '1') THEN
				IF(DW = '1') THEN
					Q <= DOUT;
				ELSE 
					Q <= D;
				END IF;
			ELSE
				Q <= Q + 1;
			END IF;
		END IF;
	END PROCESS PPC;
	
	PRAM: PROCESS(CLK) BEGIN
		IF(CLK'EVENT  AND CLK = '1') THEN
			IF(UP = '1') THEN
				STACKs(CONV_INTEGER(STACK_POINTER)) <= Q + 1;
			END IF;
		END IF;
	END PROCESS PRAM;
	
	DOUT <= STACKS(CONV_INTEGER(STACK_POINTER - 1));
end PROGRAMA;

