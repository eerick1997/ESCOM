module proyect ( 
	a,
	d
	) ;

input [1:0] a;
inout [7:0] d;
