module ffjk ( 
	j,
	k,
	clk,
	pre,
	clr,
	q,
	nq
	) ;

input  j;
input  k;
input  clk;
input  pre;
input  clr;
inout  q;
inout  nq;
