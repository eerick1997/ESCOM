module teclado ( 
	f,
	clk,
	clr,
	c,
	display
	) ;

input [3:0] f;
input  clk;
input  clr;
inout [2:0] c;
inout [6:0] display;
