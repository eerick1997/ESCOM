module ffjkyrs ( 
	j,
	k,
	clk,
	pre,
	clr,
	sel,
	q,
	nq
	) ;

input  j;
input  k;
input  clk;
input  pre;
input  clr;
input  sel;
inout  q;
inout  nq;
