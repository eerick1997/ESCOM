LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ARCHIVO_REGISTROS IS

	GENERIC(
		NBITS_ADDR : INTEGER := 4;
		NBITS_DATA : INTEGER := 16
	);
	
	PORT(
		--|============= BARREL SHIFTER =============| 
		SHAMT: IN STD_LOGIC_VECTOR( NBITS_ADDR - 1 DOWNTO 0);
		DIR : IN STD_LOGIC;		-- 1: Left Shifter , 0: Right Shifter
		
		--|=============== REGISTERS ================| 
		CLK : IN STD_LOGIC; 	--Clock
		WR : IN STD_LOGIC;	--Write Register
		
		--|======= RAM DISTRIBUTED OF 3 PORTS =======|
		ADDR_WR : IN STD_LOGIC_VECTOR( NBITS_ADDR - 1 DOWNTO 0 );	-- WRITE REGISTER
		ADDR_RD1 : IN STD_LOGIC_VECTOR( NBITS_ADDR - 1 DOWNTO 0 );	-- READ REGISTER 01
		ADDR_RD2 : IN STD_LOGIC_VECTOR( NBITS_ADDR - 1 DOWNTO 0 );	-- READ REGISTER 02
		WD : IN STD_LOGIC_VECTOR( NBITS_DATA - 1 DOWNTO 0 );		-- WRITE DATA
		DINOUT1 : INOUT STD_LOGIC_VECTOR ( NBITS_DATA - 1 DOWNTO 0);	-- READ DATA 01
		DOUT2 : OUT STD_LOGIC_VECTOR ( NBITS_DATA - 1 DOWNTO 0);	-- READ DATA 02
		SHE : IN STD_LOGIC	-- SHIFT ENABLE		
	);
	
END ARCHIVO_REGISTROS;
 
ARCHITECTURE REGISTROS OF ARCHIVO_REGISTROS IS
	
	--|=============== SIGNALS ================| 
	SIGNAL DATA_OUT : STD_LOGIC_VECTOR( NBITS_DATA - 1 DOWNTO 0 );	-- SALIDA DEL BARREL SHIFT Y ENTRADA DEL MUX
	SIGNAL DIN : STD_LOGIC_VECTOR( NBITS_DATA - 1 DOWNTO 0 );	-- DATO DE ENTRADA A LOS REGISTROS
	
	--|========== INPUT/OUTPUT FILE ===========| 
	TYPE MEM_TYPE IS ARRAY ( ( 2**NBITS_ADDR ) - 1 DOWNTO 0 ) OF STD_LOGIC_VECTOR( DIN'RANGE );
	SIGNAL MEM : MEM_TYPE;
	
	
	BEGIN
		--|======== IMPLEMENTATION OF BARREL SHIFTER ========| 
		PSHIFT : PROCESS ( SHAMT, DINOUT1, DIR )
		VARIABLE SHIFT_DATA : STD_LOGIC_VECTOR( NBITS_DATA - 1 DOWNTO 0);
		VARIABLE INDICE	: INTEGER RANGE -31 TO 32;
		
		BEGIN
			IF( DIR = '1' ) THEN 	-- 1: Left Shifter
				SHIFT_DATA := DINOUT1;
				FOR	I IN 0 TO ( NBITS_ADDR - 1 ) LOOP
					FOR J IN ( NBITS_DATA - 1 ) DOWNTO 0 LOOP
						IF( SHAMT( I ) = '1' ) THEN
							INDICE := J - 2**I;	
							IF( INDICE < 0 ) THEN	
								SHIFT_DATA( J ) := '0';
							ELSE
								SHIFT_DATA( J ) := SHIFT_DATA( INDICE );
							END IF;
						END IF;
					END LOOP;
				END LOOP;
				DATA_OUT <= SHIFT_DATA;
			ELSE						-- 0: Right Shifter
				SHIFT_DATA := DINOUT1;
				FOR	I IN 0 TO ( NBITS_ADDR - 1 ) LOOP
					FOR J IN 0 TO ( NBITS_DATA - 1 ) LOOP
						IF( SHAMT( I ) = '1' ) THEN
							INDICE := J + 2**I;	
							IF( INDICE > 7 ) THEN	
							SHIFT_DATA( J ) := '0';
							ELSE
								SHIFT_DATA( J ) := SHIFT_DATA( INDICE );
							END IF;
						END IF;
					END LOOP;
				END LOOP;
				DATA_OUT <= SHIFT_DATA;
			END IF;
		END PROCESS PSHIFT;	--CLOSE BARREL SHIFTER
		
		
		--|========== IMPLEMENTATION OF RAM DISTRIBUTED OF 3 PORTS ==========|
		
		--|================= MEMORY WRITING =================|
		PMEM : PROCESS ( CLK, SHE, WD )
		BEGIN
			-- SE ESPECIFICA EL DATO DE ESCRITURA QUE TOMA EL DATO DE ENTRADA
			IF ( SHE = '1' ) THEN
				DIN <= DATA_OUT;
			ELSE
				DIN <= WD;
			END IF;
			
			IF ( RISING_EDGE(CLK) ) THEN
				IF ( WR = '1' ) THEN 	-- WRITING
					MEM( CONV_INTEGER( ADDR_WR ) ) <= DIN;
				END IF;
			END IF;			
		END PROCESS PMEM; -- CLOSE MEMORY WRITING
		
		
		--|================= MEMORY READING =================|
		DINOUT1 <= MEM( CONV_INTEGER( ADDR_RD1 ) );
		DOUT2 <= MEM( CONV_INTEGER( ADDR_RD2 ) );
		
		-- CLOSE RAM DISTRIBUTED OF 3 PORTS
		
END REGISTROS;