library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity UNIDAD_CONTROL is
end UNIDAD_CONTROL;

architecture PROGRAMA of UNIDAD_CONTROL is

begin


end PROGRAMA;

