module det ( 
	clk,
	clr,
	e,
	s
	) ;

input  clk;
input  clr;
input  e;
inout  s;
