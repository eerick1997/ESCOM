module ffd ( 
	d,
	clk,
	pre,
	clr,
	q,
	nq
	) ;

input  d;
input  clk;
input  pre;
input  clr;
inout  q;
inout  nq;
