module dis ( 
	clr,
	clk,
	conmuta,
	display
	) ;

input  clr;
input  clk;
inout [2:0] conmuta;
inout [6:0] display;
