module ffdyt ( 
	d,
	clk,
	pre,
	clr,
	sel,
	q,
	nq
	) ;

input  d;
input  clk;
input  pre;
input  clr;
input  sel;
inout  q;
inout  nq;
