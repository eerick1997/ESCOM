module regu ( 
	clk,
	clr,
	control,
	dato,
	e
	) ;

input  clk;
input  clr;
input  control;
input [7:0] dato;
inout  e;
