module regu ( 
	clk,
	clr,
	a,
	b,
	control,
	cout,
	s0,
	s1,
	s2,
	s3,
	s4
	) ;

input  clk;
input  clr;
input  a;
input  b;
input  control;
inout  cout;
inout  s0;
inout  s1;
inout  s2;
inout  s3;
inout  s4;
