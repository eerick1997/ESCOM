module allff ( 
	clk,
	clr,
	control,
	q
	) ;

input  clk;
input  clr;
input  control;
inout [2:0] q;
