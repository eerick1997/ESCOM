library IEEE;
library work;
use IEEE.STD_LOGIC_1164.ALL;
use work.PaqueteEscomips.all;

ENTITY PROCESADOR IS
	PORT ( 
		CLK	: IN STD_LOGIC;
		CLR	: IN STD_LOGIC;
		DATAIN : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) -- SALIDA DE LA ALU
		--ADDRESS	: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		--WD : OUT STD_LOGIC
	);
END PROCESADOR;

ARCHITECTURE Behavioral OF PROCESADOR IS

SIGNAL INS					:  STD_LOGIC_VECTOR(19 DOWNTO 0);

	--INS(19) = UP
	--INS(18) = DW
	--INS(17) = WPC
	--INS(16) = SDMP
	--INS(15) = SR2
	--INS(14) = SWD
	--INS(13) = SHE
	--INS(12) = DIR
	--INS(11) = WR
	--INS(10) = LF
	--INS(9)  = SEXT
	--INS(8)  = SOP1
	--INS(7)  = SOP2
	--INS(6:3)= ALUOP
	--INS(2)  = SDMD
	--INS(1)  = WD
	--INS(0)  = SR

-- OSCILADOR DE DIVISOR DE FRECUENCIA
SIGNAL OSC					: STD_LOGIC;

-- BUSES
SIGNAL BUS_AZUL			:	STD_LOGIC_VECTOR(15 DOWNTO 0); -- PILA -> MEMORIA DE PROGRAMA && SOP1
SIGNAL BUS_NEGRO			:  STD_LOGIC_VECTOR(24 DOWNTO 0);

-- SALIDAS DE LOS MUXES
SIGNAL MUX_SR2				:	STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL MUX_SWD				:	STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MUX_SDMP			:	STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MUX_SEXT			:	STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MUX_SOP1			:	STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MUX_SOP2			:	STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MUX_SDMD			:  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL MUX_SR				:  STD_LOGIC_VECTOR(15 DOWNTO 0);

-- SALIDAS ARCHIVO DE REGISTRO
SIGNAL READ_DATA1			:	STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL READ_DATA2			:	STD_LOGIC_VECTOR(15 DOWNTO 0);

-- SALIDAS EXTENSORES
SIGNAL EXTENSOR_SIGNO	:	STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL EXTENSOR_DIREC	:	STD_LOGIC_VECTOR(15 DOWNTO 0);

--- SALIDAS MEMORIA DE DATOS
SIGNAL MEMORIA_DATOS_D	:	STD_LOGIC_VECTOR(15 DOWNTO 0);

-- SALIDAS ALU
SIGNAL ALU_D				:	STD_LOGIC_VECTOR(15 DOWNTO 0);	

-- ENTRADAS PILA
SIGNAL PILA_D				:  STD_LOGIC_VECTOR(15 DOWNTO 0);

-- ENTRADAS MEMORIA DE PROGRAMA
SIGNAL MEMORIA_PROG_A	:	STD_LOGIC_VECTOR(15 DOWNTO 0);

-- ENTRADAS ARCHIVO DE REGISTRO
SIGNAL READ_REGISTER1	:	STD_LOGIC_VECTOR(3 DOWNTO 0);

-- SALIDAS DE CONTROL
SIGNAL BANDERAS			:  STD_LOGIC_VECTOR(3 DOWNTO 0);
-- PILA

BEGIN

--	DIV	: DIVISOR PORT MAP(
--		OSC_CLK		=> 	OSC_CLK,
--		CLR			=>	CLR,
--		CLK			=>	CLK
--	);

	FREC: DIVISOR_FRECUENCIA PORT MAP(
		OSC=>CLK,
		CLR=>CLR,
		CLK=>OSC
	);	
	
	MEM_PROGRAMA: MEMORIA_PROGRAMA PORT MAP(
		A => BUS_AZUL,
		D => BUS_NEGRO
	);
	
	STACK: PILA PORT MAP(
		CLK => OSC,
		CLR => CLR,
		WPC => INS(17),
		UP	 => INS(19),
		DW  => INS(18),
		D   => MUX_SDMP,
		Q   => BUS_AZUL
	);
	
	PRIN_CONTROL: PRINCIPAL_CONTROL PORT MAP(
		CLK		=>	OSC,
		CLR		=> CLR,
		LF			=> INS(10),	
		MICRO		=> INS,
		FUNCODE 	=> BUS_NEGRO(3 DOWNTO 0),
		OPCODE	=> BUS_NEGRO(24 DOWNTO 20),
		BANDERAS => BANDERAS
	);
	
	ARCH_REGISTROS: ARCHIVO_REGISTROS PORT MAP(
		CLK 		=>	OSC,
		SHAMT 	=> BUS_NEGRO(7 DOWNTO 4),
		DIR 		=> INS(12),
		WR 		=> INS(11), 
		ADDR_WR 	=> BUS_NEGRO(19 DOWNTO 16),
		ADDR_RD1 => BUS_NEGRO(15 DOWNTO 12),
		ADDR_RD2 => MUX_SR2,
		WD			=> MUX_SWD,
		DINOUT1  => READ_DATA1,
		DOUT2		=> READ_DATA2,
		SHE		=> INS(13)
	);
	
	UAL: ALU PORT MAP(
		A 			=> MUX_SOP1,
		B			=> MUX_SOP2,
		ALUOP		=> INS(6 DOWNTO 3),
		RES		=> ALU_D,
		FLAGS		=> BANDERAS
	);
	
	MEM_DATOS: MEMORIA_DATOS PORT MAP(
		CLK 					=>	OSC,
		BUS_DATOS_ENTRADA =>	READ_DATA2,
		BUS_DATOS_SALIDA  => MEMORIA_DATOS_D,
		ADR					=> MUX_SDMD,
		WD						=> INS(1)	
	);
	
	MUX_SR <= ALU_D WHEN (INS(0) = '1') ELSE MEMORIA_DATOS_D;
	
	EXTENSOR_SIGNO <= X"F"&BUS_NEGRO(11 DOWNTO 0) WHEN(BUS_NEGRO(11) = '1')
					 ELSE X"0"&BUS_NEGRO(11 DOWNTO 0);

	EXTENSOR_DIREC <= X"0"&BUS_NEGRO(11 DOWNTO 0);
	
	MUX_SDMP <= MUX_SR WHEN INS(16) = '1' ELSE BUS_NEGRO( 15 DOWNTO 0);
	MUX_SEXT <= EXTENSOR_DIREC WHEN INS(9) = '1' ELSE EXTENSOR_SIGNO;
	
	MUX_SWD  <= MUX_SR WHEN INS(14) = '1' ELSE BUS_NEGRO (15 DOWNTO 0);
	MUX_SR2  <= BUS_NEGRO (19 DOWNTO 16) WHEN INS(15) = '1' ELSE 
					BUS_NEGRO (11 DOWNTO 8 );
	
	MUX_SOP1 <= BUS_AZUL WHEN (INS(8) = '1') ELSE READ_DATA1;
	MUX_SOP2 <= MUX_SEXT WHEN (INS(7) = '1') ELSE READ_DATA2;
	
	MUX_SDMD <= BUS_NEGRO(15 DOWNTO 0) WHEN (INS(2) = '1') ELSE ALU_D;
	
	DATAIN 	<= 	READ_DATA2;
	
END Behavioral;

