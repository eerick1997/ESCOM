module regu ( 
	clk,
	clr,
	control,
	dato1,
	dato2,
	a,
	b
	) ;

input  clk;
input  clr;
input  control;
input [3:0] dato1;
input [3:0] dato2;
inout  a;
inout  b;
