module p11 ( 
	clk,
	clr,
	change,
	display
	) ;

input  clk;
input  clr;
inout [2:0] change;
inout [6:0] display;
